LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
ENTITY lights IS
PORT (
SW : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
KEY : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
CLOCK_50 : IN STD_LOGIC;
DRAM_CLK, DRAM_CKE : OUT STD_LOGIC;
LEDG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
DRAM_ADDR : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
DRAM_BA_1, DRAM_BA_0 : BUFFER STD_LOGIC;
DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N, DRAM_WE_N : OUT STD_LOGIC;
DRAM_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
DRAM_UDQM, DRAM_LDQM : BUFFER STD_LOGIC
);
END lights;

ARCHITECTURE Structure OF lights IS
COMPONENT nios_system
PORT (
clk_0 : IN STD_LOGIC;
reset_n : IN STD_LOGIC;
out_port_from_the_LED_S : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
in_port_to_the_Switches : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
zs_addr_from_the_sdram_1: OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
zs_ba_from_the_sdram_1: BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0);
zs_cas_n_from_the_sdram_1: OUT STD_LOGIC;
zs_cke_from_the_sdram_1: OUT STD_LOGIC;
zs_cs_n_from_the_sdram_1: OUT STD_LOGIC;
zs_dq_to_and_from_the_sdram_1: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
zs_dqm_from_the_sdram_1: BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0);
zs_ras_n_from_the_sdram_1: OUT STD_LOGIC;
zs_we_n_from_the_sdram_1: OUT STD_LOGIC );
END COMPONENT;
COMPONENT sdram_1_pll
PORT ( inclk0 : IN STD_LOGIC;
c0 : OUT STD_LOGIC );
END COMPONENT;
SIGNAL BA : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL DQM : STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
BA <= (DRAM_BA_1 & DRAM_BA_0);
DQM <= (DRAM_UDQM & DRAM_LDQM);
-- Instantiate the Nios II system entity generated by the SOPC Builder
NiosII: nios_system PORT MAP (CLOCK_50, KEY(0), LEDG, SW,
DRAM_ADDR, BA, DRAM_CAS_N, DRAM_CKE, DRAM_CS_N,
DRAM_DQ, DQM, DRAM_RAS_N, DRAM_WE_N );
DRAM_CLK <= CLOCK_50;
END Structure;